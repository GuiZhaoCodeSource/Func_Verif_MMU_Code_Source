/******************************************************************************
* (C) Copyright 2011 KALRAY SA All Rights Reserved
*
* MODULE:    mmucfg.svh
* DEVICE:    MMUCFG VIP
* PROJECT:
* AUTHOR:
* DATE:
*
* ABSTRACT:
*
*******************************************************************************/
`ifndef MMUCFG_SVH
`define MMUCFG_SVH

// Include
`include "mmucfg_transfer.sv"
`include "mmucfg_master_sequencer.sv"
`include "mmucfg_master_driver.sv"
`include "mmucfg_master_agent.sv"
`include "mmucfg_slave_sequencer.sv"
`include "mmucfg_slave_driver.sv"
`include "mmucfg_slave_agent.sv"
`include "mmucfg_bus_monitor.sv"
`include "mmucfg_env.sv"
`endif
