/******************************************************************************
* (C) Copyright 2011 KALRAY SA All Rights Reserved
*
* MODULE:    mmu_proc_tlbmaintenance.svh
* DEVICE:    MMU_PROC_TLBMAINTENANCE VIP
* PROJECT:
* AUTHOR:
* DATE:
*
* ABSTRACT:
*
*******************************************************************************/
`ifndef MMU_PROC_TLBMAINTENANCE_SVH
`define MMU_PROC_TLBMAINTENANCE_SVH

// Include
`include "mmu_proc_tlbmaintenance_transfer.sv"
`include "mmu_proc_tlbmaintenance_master_sequencer.sv"
`include "mmu_proc_tlbmaintenance_master_driver.sv"
`include "mmu_proc_tlbmaintenance_master_agent.sv"
`include "mmu_proc_tlbmaintenance_slave_sequencer.sv"
`include "mmu_proc_tlbmaintenance_slave_driver.sv"
`include "mmu_proc_tlbmaintenance_slave_agent.sv"
`include "mmu_proc_tlbmaintenance_bus_monitor.sv"
`include "mmu_proc_tlbmaintenance_env.sv"
`endif
